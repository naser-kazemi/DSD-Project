module rope (

);

endmodule