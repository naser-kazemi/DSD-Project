module FixPointALU (
    input wire[31:0] in_1,
);
    
endmodule