`include "FixedPointALU.v"


module EnforceConstraints (
    input wire[31:0] up_x_pos,
    input wire[31:0] up_y_pos,
    input wire[31:0] x_pos,
    input wire[31:0] y_pos,
    input wire[31:0] down_x_pos,
    input wire[31:0] down_y_pos,
    output [31:0] x_enforced_constraints,
    output [31:0] y_enforced_constraints
);









endmodule